`timescale 1ns / 1ps
/*************************************************************************************
    Mealy型电路两段式独热码检测比特流序列10101011
    输入：x(单个比特数字)、rstn(低电平有效状态清零)、clk(时钟信号，每次输入产生一个时钟信号)；
    输出：y(是否存在序列，若出现序列则不计算前面重叠部分)、s(8位独热码led显示当前状态)。
*************************************************************************************/
module FSM2(
    input x,rstn,clk,
    output reg y,
    output reg[7:0] s
);
    reg[7:0] d,q;//s的次态与现态
    reg y_ns,y_cs;//y的次态与现态
    always @(*)begin//通过现态与输入计算次态
        d[7]=q[6]&&x;
        d[6]=q[5]&&(~x);
        d[5]=q[4]&&x;
        d[4]=q[3]&&(~x);
        d[3]=q[2]&&x;
        d[2]=q[1]&&(~x);
        d[1]=x&&(q[0]||q[1]||q[3]||q[5]);
        d[0]=(x&&q[7])||((~x)&&(q[0]||q[2]||q[4]||q[6]||q[7]));       
        y_ns=q[7]&&x;
        y=y_cs;
        s=q;
    end
    always @(posedge clk , negedge rstn)
    begin
        if(!rstn)begin//接收到清零信号
            q[7:0]<=8'h01;
        end
        else begin//更新状态
            y_cs<=y_ns;
            q[7:0]<=d[7:0];
        end
    end
endmodule